##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri May 27 22:50:21 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 829.380000 BY 820.080000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.3816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.976 LAYER met3  ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 15.1 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.311 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1.625000 0.000000 1.765000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.6426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.987 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 37.839 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 187.983 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 9.960000 0.490000 10.100000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.315000 0.000000 176.455000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.290000 0.000000 59.430000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.010000 0.000000 178.150000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.620000 0.000000 174.760000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.920000 0.000000 173.060000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.225000 0.000000 171.365000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.530000 0.000000 169.670000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.560000 0.000000 113.700000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.865000 0.000000 112.005000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.170000 0.000000 110.310000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.475000 0.000000 108.615000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.780000 0.000000 106.920000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.080000 0.000000 105.220000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.385000 0.000000 103.525000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.690000 0.000000 101.830000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.995000 0.000000 100.135000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.300000 0.000000 98.440000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.600000 0.000000 96.740000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.905000 0.000000 95.045000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.210000 0.000000 93.350000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.515000 0.000000 91.655000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.820000 0.000000 89.960000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.120000 0.000000 88.260000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.425000 0.000000 86.565000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730000 0.000000 84.870000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.035000 0.000000 83.175000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.340000 0.000000 81.480000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.640000 0.000000 79.780000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.945000 0.000000 78.085000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.250000 0.000000 76.390000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.555000 0.000000 74.695000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.860000 0.000000 73.000000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.160000 0.000000 71.300000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.465000 0.000000 69.605000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.770000 0.000000 67.910000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.075000 0.000000 66.215000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.380000 0.000000 64.520000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.680000 0.000000 62.820000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.985000 0.000000 61.125000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.595000 0.000000 57.735000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.900000 0.000000 56.040000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.200000 0.000000 54.340000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.505000 0.000000 52.645000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.810000 0.000000 50.950000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.115000 0.000000 49.255000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.420000 0.000000 47.560000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.720000 0.000000 45.860000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.025000 0.000000 44.165000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.330000 0.000000 42.470000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.635000 0.000000 40.775000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.940000 0.000000 39.080000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.240000 0.000000 37.380000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.545000 0.000000 35.685000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.850000 0.000000 33.990000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.155000 0.000000 32.295000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.460000 0.000000 30.600000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.760000 0.000000 28.900000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.065000 0.000000 27.205000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.370000 0.000000 25.510000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.675000 0.000000 23.815000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.980000 0.000000 22.120000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.280000 0.000000 20.420000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.585000 0.000000 18.725000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.890000 0.000000 17.030000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.195000 0.000000 15.335000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.500000 0.000000 13.640000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.800000 0.000000 11.940000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.105000 0.000000 10.245000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.410000 0.000000 8.550000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.715000 0.000000 6.855000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.020000 0.000000 5.160000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.651 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 3.320000 0.000000 3.460000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.031 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 167.835000 0.000000 167.975000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 166.140000 0.000000 166.280000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.440000 0.000000 164.580000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.745000 0.000000 162.885000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 161.050000 0.000000 161.190000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 159.355000 0.000000 159.495000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 157.660000 0.000000 157.800000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.960000 0.000000 156.100000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 154.265000 0.000000 154.405000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 152.570000 0.000000 152.710000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 150.875000 0.000000 151.015000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 149.180000 0.000000 149.320000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 147.480000 0.000000 147.620000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 145.785000 0.000000 145.925000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 144.090000 0.000000 144.230000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 142.395000 0.000000 142.535000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 140.700000 0.000000 140.840000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 139.000000 0.000000 139.140000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 137.305000 0.000000 137.445000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 135.610000 0.000000 135.750000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 133.915000 0.000000 134.055000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 132.220000 0.000000 132.360000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 130.520000 0.000000 130.660000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 128.825000 0.000000 128.965000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 127.130000 0.000000 127.270000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 125.435000 0.000000 125.575000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 123.740000 0.000000 123.880000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 122.040000 0.000000 122.180000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 120.345000 0.000000 120.485000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 118.650000 0.000000 118.790000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.08 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 116.955000 0.000000 117.095000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.884 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 115.260000 0.000000 115.400000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.100000 0.000000 395.240000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.400000 0.000000 393.540000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.705000 0.000000 391.845000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.010000 0.000000 390.150000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.315000 0.000000 388.455000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.620000 0.000000 386.760000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.920000 0.000000 385.060000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.225000 0.000000 383.365000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.530000 0.000000 381.670000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.835000 0.000000 379.975000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.140000 0.000000 378.280000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.440000 0.000000 376.580000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.745000 0.000000 374.885000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.050000 0.000000 373.190000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.355000 0.000000 371.495000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.660000 0.000000 369.800000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.960000 0.000000 368.100000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.265000 0.000000 366.405000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.570000 0.000000 364.710000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.875000 0.000000 363.015000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.180000 0.000000 361.320000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.480000 0.000000 359.620000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.785000 0.000000 357.925000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.090000 0.000000 356.230000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.395000 0.000000 354.535000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.700000 0.000000 352.840000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.000000 0.000000 351.140000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.305000 0.000000 349.445000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.610000 0.000000 347.750000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.915000 0.000000 346.055000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.220000 0.000000 344.360000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.520000 0.000000 342.660000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.825000 0.000000 340.965000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.130000 0.000000 339.270000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.435000 0.000000 337.575000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.740000 0.000000 335.880000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.040000 0.000000 334.180000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.345000 0.000000 332.485000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.650000 0.000000 330.790000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.955000 0.000000 329.095000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.260000 0.000000 327.400000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.560000 0.000000 325.700000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.865000 0.000000 324.005000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.170000 0.000000 322.310000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.475000 0.000000 320.615000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.780000 0.000000 318.920000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.080000 0.000000 317.220000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.385000 0.000000 315.525000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.690000 0.000000 313.830000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.995000 0.000000 312.135000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.300000 0.000000 310.440000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.600000 0.000000 308.740000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.905000 0.000000 307.045000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.210000 0.000000 305.350000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.515000 0.000000 303.655000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.820000 0.000000 301.960000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.120000 0.000000 300.260000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.425000 0.000000 298.565000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.730000 0.000000 296.870000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.035000 0.000000 295.175000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.340000 0.000000 293.480000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.640000 0.000000 291.780000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.87 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 234.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 64.5348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 344.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2075 LAYER met4  ;
    ANTENNAMAXAREACAR 17.5775 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 92.0002 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.22669 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 289.945000 0.000000 290.085000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 234.286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1254.69 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 10.125 LAYER met4  ;
    ANTENNAMAXAREACAR 83.8539 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 427.107 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.662917 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 288.250000 0.000000 288.390000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.555000 0.000000 286.695000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.860000 0.000000 285.000000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.160000 0.000000 283.300000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.465000 0.000000 281.605000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770000 0.000000 279.910000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.075000 0.000000 278.215000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.380000 0.000000 276.520000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.680000 0.000000 274.820000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.985000 0.000000 273.125000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.290000 0.000000 271.430000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.595000 0.000000 269.735000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.900000 0.000000 268.040000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.200000 0.000000 266.340000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.505000 0.000000 264.645000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.810000 0.000000 262.950000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.115000 0.000000 261.255000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.420000 0.000000 259.560000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.720000 0.000000 257.860000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.025000 0.000000 256.165000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.330000 0.000000 254.470000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.635000 0.000000 252.775000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.940000 0.000000 251.080000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.240000 0.000000 249.380000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.545000 0.000000 247.685000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.850000 0.000000 245.990000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.155000 0.000000 244.295000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.460000 0.000000 242.600000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.760000 0.000000 240.900000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.065000 0.000000 239.205000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.370000 0.000000 237.510000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.675000 0.000000 235.815000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.980000 0.000000 234.120000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.280000 0.000000 232.420000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.585000 0.000000 230.725000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.890000 0.000000 229.030000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.195000 0.000000 227.335000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.500000 0.000000 225.640000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.800000 0.000000 223.940000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.105000 0.000000 222.245000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.410000 0.000000 220.550000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.715000 0.000000 218.855000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.020000 0.000000 217.160000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.320000 0.000000 215.460000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.625000 0.000000 213.765000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.930000 0.000000 212.070000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.235000 0.000000 210.375000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.540000 0.000000 208.680000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.840000 0.000000 206.980000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.145000 0.000000 205.285000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.450000 0.000000 203.590000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.755000 0.000000 201.895000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.060000 0.000000 200.200000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.360000 0.000000 198.500000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.665000 0.000000 196.805000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.970000 0.000000 195.110000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.275000 0.000000 193.415000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.580000 0.000000 191.720000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.880000 0.000000 190.020000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.185000 0.000000 188.325000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.490000 0.000000 186.630000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.795000 0.000000 184.935000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.100000 0.000000 183.240000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7324 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.6195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 181.400000 0.000000 181.540000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.705000 0.000000 179.845000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 612.185000 0.000000 612.325000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 610.490000 0.000000 610.630000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 608.795000 0.000000 608.935000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 607.100000 0.000000 607.240000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 605.400000 0.000000 605.540000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 603.705000 0.000000 603.845000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 602.010000 0.000000 602.150000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 600.315000 0.000000 600.455000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 598.620000 0.000000 598.760000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 596.920000 0.000000 597.060000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 595.225000 0.000000 595.365000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 593.530000 0.000000 593.670000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 591.835000 0.000000 591.975000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 590.140000 0.000000 590.280000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 588.440000 0.000000 588.580000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 586.745000 0.000000 586.885000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 585.050000 0.000000 585.190000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 583.355000 0.000000 583.495000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 581.660000 0.000000 581.800000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 579.960000 0.000000 580.100000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 578.265000 0.000000 578.405000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 576.570000 0.000000 576.710000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 574.875000 0.000000 575.015000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 573.180000 0.000000 573.320000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 571.480000 0.000000 571.620000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 569.785000 0.000000 569.925000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 568.090000 0.000000 568.230000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 566.395000 0.000000 566.535000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 564.700000 0.000000 564.840000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 563.000000 0.000000 563.140000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 561.305000 0.000000 561.445000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 559.610000 0.000000 559.750000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 557.915000 0.000000 558.055000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 556.220000 0.000000 556.360000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 554.520000 0.000000 554.660000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 552.825000 0.000000 552.965000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 551.130000 0.000000 551.270000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 549.435000 0.000000 549.575000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 547.740000 0.000000 547.880000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 546.040000 0.000000 546.180000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 544.345000 0.000000 544.485000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 542.650000 0.000000 542.790000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 540.955000 0.000000 541.095000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 539.260000 0.000000 539.400000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 537.560000 0.000000 537.700000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 535.865000 0.000000 536.005000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 534.170000 0.000000 534.310000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 532.475000 0.000000 532.615000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 530.780000 0.000000 530.920000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 529.080000 0.000000 529.220000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 527.385000 0.000000 527.525000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 525.690000 0.000000 525.830000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 523.995000 0.000000 524.135000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 522.300000 0.000000 522.440000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 520.600000 0.000000 520.740000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 518.905000 0.000000 519.045000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 517.210000 0.000000 517.350000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 515.515000 0.000000 515.655000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 513.820000 0.000000 513.960000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 512.120000 0.000000 512.260000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 510.425000 0.000000 510.565000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 508.730000 0.000000 508.870000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 507.035000 0.000000 507.175000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 505.340000 0.000000 505.480000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 503.640000 0.000000 503.780000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.613 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 501.945000 0.000000 502.085000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 500.250000 0.000000 500.390000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 498.555000 0.000000 498.695000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 496.860000 0.000000 497.000000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 495.160000 0.000000 495.300000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 493.465000 0.000000 493.605000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 491.770000 0.000000 491.910000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 490.075000 0.000000 490.215000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 488.380000 0.000000 488.520000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 486.680000 0.000000 486.820000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 484.985000 0.000000 485.125000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 483.290000 0.000000 483.430000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 481.595000 0.000000 481.735000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 479.900000 0.000000 480.040000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 478.200000 0.000000 478.340000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 476.505000 0.000000 476.645000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 474.810000 0.000000 474.950000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 473.115000 0.000000 473.255000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 471.420000 0.000000 471.560000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 469.720000 0.000000 469.860000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 468.025000 0.000000 468.165000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 466.330000 0.000000 466.470000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 464.635000 0.000000 464.775000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 462.940000 0.000000 463.080000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 461.240000 0.000000 461.380000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 459.545000 0.000000 459.685000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 457.850000 0.000000 457.990000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 456.155000 0.000000 456.295000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 454.460000 0.000000 454.600000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 452.760000 0.000000 452.900000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 451.065000 0.000000 451.205000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 449.370000 0.000000 449.510000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 447.675000 0.000000 447.815000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 445.980000 0.000000 446.120000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 444.280000 0.000000 444.420000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 442.585000 0.000000 442.725000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.253 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 440.890000 0.000000 441.030000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 439.195000 0.000000 439.335000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.554 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 437.500000 0.000000 437.640000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.98 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 435.800000 0.000000 435.940000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.456 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 434.105000 0.000000 434.245000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.79 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 432.410000 0.000000 432.550000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 430.715000 0.000000 430.855000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.05 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 429.020000 0.000000 429.160000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.84 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 427.320000 0.000000 427.460000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.578 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 425.625000 0.000000 425.765000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.307 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 423.930000 0.000000 424.070000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 422.235000 0.000000 422.375000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 420.540000 0.000000 420.680000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 418.840000 0.000000 418.980000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 417.145000 0.000000 417.285000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 415.450000 0.000000 415.590000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 413.755000 0.000000 413.895000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 412.060000 0.000000 412.200000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 410.360000 0.000000 410.500000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 408.665000 0.000000 408.805000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 406.970000 0.000000 407.110000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 405.275000 0.000000 405.415000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 403.580000 0.000000 403.720000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 401.880000 0.000000 402.020000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 400.185000 0.000000 400.325000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 398.490000 0.000000 398.630000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.242 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 396.795000 0.000000 396.935000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.500000 0.000000 818.640000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.580000 0.000000 827.720000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.880000 0.000000 826.020000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.185000 0.000000 824.325000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.490000 0.000000 822.630000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.795000 0.000000 820.935000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.100000 0.000000 819.240000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.400000 0.000000 817.540000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.705000 0.000000 815.845000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.010000 0.000000 814.150000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.315000 0.000000 812.455000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.620000 0.000000 810.760000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.920000 0.000000 809.060000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.225000 0.000000 807.365000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.530000 0.000000 805.670000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.835000 0.000000 803.975000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.140000 0.000000 802.280000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.440000 0.000000 800.580000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.745000 0.000000 798.885000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.050000 0.000000 797.190000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.355000 0.000000 795.495000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.660000 0.000000 793.800000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.960000 0.000000 792.100000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.265000 0.000000 790.405000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.570000 0.000000 788.710000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.875000 0.000000 787.015000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.180000 0.000000 785.320000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.480000 0.000000 783.620000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.785000 0.000000 781.925000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.090000 0.000000 780.230000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.395000 0.000000 778.535000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.700000 0.000000 776.840000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.000000 0.000000 775.140000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.305000 0.000000 773.445000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.610000 0.000000 771.750000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.915000 0.000000 770.055000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.220000 0.000000 768.360000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.520000 0.000000 766.660000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.825000 0.000000 764.965000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.130000 0.000000 763.270000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.435000 0.000000 761.575000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.740000 0.000000 759.880000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.040000 0.000000 758.180000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.345000 0.000000 756.485000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.650000 0.000000 754.790000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.955000 0.000000 753.095000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.260000 0.000000 751.400000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.560000 0.000000 749.700000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.865000 0.000000 748.005000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.170000 0.000000 746.310000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.475000 0.000000 744.615000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.780000 0.000000 742.920000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.080000 0.000000 741.220000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.385000 0.000000 739.525000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.690000 0.000000 737.830000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.995000 0.000000 736.135000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.300000 0.000000 734.440000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.600000 0.000000 732.740000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.905000 0.000000 731.045000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.210000 0.000000 729.350000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.515000 0.000000 727.655000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.820000 0.000000 725.960000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 78.163 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 417.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 59.6178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.92 LAYER met4  ;
    ANTENNAMAXAREACAR 8.69213 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 45.2602 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0474242 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 724.120000 0.000000 724.260000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 137.414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 735.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 15.36 LAYER met4  ;
    ANTENNAMAXAREACAR 59.9743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 313.116 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.357563 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 722.425000 0.000000 722.565000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.730000 0.000000 720.870000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.035000 0.000000 719.175000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.340000 0.000000 717.480000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.640000 0.000000 715.780000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.945000 0.000000 714.085000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.250000 0.000000 712.390000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.555000 0.000000 710.695000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.860000 0.000000 709.000000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.160000 0.000000 707.300000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.465000 0.000000 705.605000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.770000 0.000000 703.910000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.075000 0.000000 702.215000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.380000 0.000000 700.520000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.680000 0.000000 698.820000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.985000 0.000000 697.125000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.290000 0.000000 695.430000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.595000 0.000000 693.735000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.900000 0.000000 692.040000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.200000 0.000000 690.340000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.505000 0.000000 688.645000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.810000 0.000000 686.950000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.115000 0.000000 685.255000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.420000 0.000000 683.560000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.720000 0.000000 681.860000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.025000 0.000000 680.165000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.330000 0.000000 678.470000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.635000 0.000000 676.775000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.940000 0.000000 675.080000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.240000 0.000000 673.380000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.545000 0.000000 671.685000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850000 0.000000 669.990000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.155000 0.000000 668.295000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.994 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.1503 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 666.460000 0.000000 666.600000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.302 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.83232 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.1253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 664.760000 0.000000 664.900000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.95253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.6101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 663.065000 0.000000 663.205000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.729 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2866 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.2667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 661.370000 0.000000 661.510000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.25131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.5394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 659.675000 0.000000 659.815000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.134 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.21737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.0545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 657.980000 0.000000 658.120000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.316 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.54667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.9939 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 656.280000 0.000000 656.420000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.03 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 654.585000 0.000000 654.725000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.833 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.76 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.5374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 652.890000 0.000000 653.030000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.42222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.0747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 651.195000 0.000000 651.335000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.533 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.57636 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.7293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 649.500000 0.000000 649.640000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.554 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.69707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.1152 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 647.800000 0.000000 647.940000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.554 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.96667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4768 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 646.105000 0.000000 646.245000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.34717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.8424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 644.410000 0.000000 644.550000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.9841 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 642.715000 0.000000 642.855000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2278 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.6111 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 641.020000 0.000000 641.160000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.320000 0.000000 639.460000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.625000 0.000000 637.765000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.930000 0.000000 636.070000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.235000 0.000000 634.375000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.540000 0.000000 632.680000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.840000 0.000000 630.980000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.145000 0.000000 629.285000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.450000 0.000000 627.590000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.755000 0.000000 625.895000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.060000 0.000000 624.200000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.360000 0.000000 622.500000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.665000 0.000000 620.805000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.970000 0.000000 619.110000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.275000 0.000000 617.415000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.973 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.2563 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.161635 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 615.580000 0.000000 615.720000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.880000 0.000000 614.020000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.850000 0.800000 40.150000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 99.855000 0.800000 100.155000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 159.860000 0.800000 160.160000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 219.860000 0.800000 220.160000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 279.865000 0.800000 280.165000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 339.865000 0.800000 340.165000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 399.870000 0.800000 400.170000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 459.875000 0.800000 460.175000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 519.875000 0.800000 520.175000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 579.880000 0.800000 580.180000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 639.880000 0.800000 640.180000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 699.885000 0.800000 700.185000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 759.890000 0.800000 760.190000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.830000 0.800000 11.130000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.730000 819.590000 63.870000 820.080000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.425000 819.590000 159.565000 820.080000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.120000 819.590000 255.260000 820.080000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.820000 819.590000 350.960000 820.080000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.515000 819.590000 446.655000 820.080000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.215000 819.590000 542.355000 820.080000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.910000 819.590000 638.050000 820.080000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.605000 819.590000 733.745000 820.080000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.880000 819.590000 820.020000 820.080000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 782.645000 829.380000 782.945000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 726.730000 829.380000 727.030000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 670.820000 829.380000 671.120000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 614.905000 829.380000 615.205000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 558.990000 829.380000 559.290000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 503.075000 829.380000 503.375000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 447.160000 829.380000 447.460000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 391.250000 829.380000 391.550000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 335.335000 829.380000 335.635000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 124.4 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 645.641 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 12.9226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.912 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 13.0528 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.1887 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 279.420000 829.380000 279.720000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 223.505000 829.380000 223.805000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 167.590000 829.380000 167.890000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 111.680000 829.380000 111.980000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 55.765000 829.380000 56.065000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 828.580000 9.610000 829.380000 9.910000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.850000 0.800000 20.150000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.855000 0.800000 80.155000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 139.855000 0.800000 140.155000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 199.860000 0.800000 200.160000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 259.865000 0.800000 260.165000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 319.865000 0.800000 320.165000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 379.870000 0.800000 380.170000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 439.870000 0.800000 440.170000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.221 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.62 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 499.875000 0.800000 500.175000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 559.880000 0.800000 560.180000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 619.880000 0.800000 620.180000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 679.885000 0.800000 680.185000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 739.885000 0.800000 740.185000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 799.890000 0.800000 800.190000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 431.661 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2275.67 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.2064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 186.382 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 994.976 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 1490.14 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 7949.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 31.830000 819.590000 31.970000 820.080000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5628 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.653 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8591 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.6746 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.4224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 262.016 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 389.819 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2101.58 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 186.176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 993.872 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 1485.12 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 7924.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 127.525000 819.590000 127.665000 820.080000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 361.672 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1922.87 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.0938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 186.111 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 994 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 1529.67 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 8152.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 223.225000 819.590000 223.365000 820.080000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 208.427 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1113.02 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 1694.73 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 9035.52 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 8.6889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.1655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.7174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.904 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 373.391 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1974.56 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 318.920000 819.590000 319.060000 820.080000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 335.125 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1780.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 27.1918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.562 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.232 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.704 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 403.882 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2144.36 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 414.615000 819.590000 414.755000 820.080000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 66.0849 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 351.611 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 66.4453 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 331.594 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.5999 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 211.664 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 429.318 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2279.33 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 510.315000 819.590000 510.455000 820.080000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 21.7607 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.4167 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 23.752 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.766 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.1165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.831 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 323.824 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 511.286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2731.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 606.010000 819.590000 606.150000 820.080000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.6837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.115 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 33.3107 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.829 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.1623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.533 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7357 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.1792 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.504 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 504.592 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2669.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 701.710000 819.590000 701.850000 820.080000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 98.5618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 528.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 98.9944 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 528.373 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 797.405000 819.590000 797.545000 820.080000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 94.2961 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 505.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 128.331 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 666.96 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 801.285000 829.380000 801.585000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 89.9369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 476.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 105.047 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 561.52 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 285.544 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1513.29 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 745.370000 829.380000 745.670000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 101.011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 542.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 75.7643 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.294 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 689.455000 829.380000 689.755000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 110.124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 590.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 123.258 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 646.127 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 633.540000 829.380000 633.840000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.8546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 513.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 177.76 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 938.563 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 577.630000 829.380000 577.930000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.5617 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 301.676 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1613.76 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 521.715000 829.380000 522.015000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.3882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 196.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 331.606 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1770.63 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.2846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 471.792 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 707.832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3778.93 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 465.800000 829.380000 466.100000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 409.885000 829.380000 410.185000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.78 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 353.970000 829.380000 354.270000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 298.060000 829.380000 298.360000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 242.145000 829.380000 242.445000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 186.230000 829.380000 186.530000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 130.315000 829.380000 130.615000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 74.400000 829.380000 74.700000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 18.490000 829.380000 18.790000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.221 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.95 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 10.200000 0.000000 10.500000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.855000 0.800000 60.155000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.855000 0.800000 120.155000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 179.860000 0.800000 180.160000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 239.860000 0.800000 240.160000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 299.865000 0.800000 300.165000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 359.870000 0.800000 360.170000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 419.870000 0.800000 420.170000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 479.875000 0.800000 480.175000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 539.875000 0.800000 540.175000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 599.880000 0.800000 600.180000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 659.885000 0.800000 660.185000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 719.885000 0.800000 720.185000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 779.890000 0.800000 780.190000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 10.280000 819.590000 10.420000 820.080000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 95.625000 819.590000 95.765000 820.080000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 191.325000 819.590000 191.465000 820.080000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 287.020000 819.590000 287.160000 820.080000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.456 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 382.720000 819.590000 382.860000 820.080000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 478.415000 819.590000 478.555000 820.080000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 574.110000 819.590000 574.250000 820.080000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 669.810000 819.590000 669.950000 820.080000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 379.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 765.505000 819.590000 765.645000 820.080000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.78 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 819.690000 829.380000 819.990000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 764.010000 829.380000 764.310000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 708.095000 829.380000 708.395000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 652.180000 829.380000 652.480000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 596.265000 829.380000 596.565000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 540.350000 829.380000 540.650000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 484.440000 829.380000 484.740000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 428.525000 829.380000 428.825000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.78 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 372.610000 829.380000 372.910000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 122.915 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 656.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 64.9637 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 349.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.156 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5704 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.928175 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 316.695000 829.380000 316.995000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 260.780000 829.380000 261.080000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 204.870000 829.380000 205.170000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 148.955000 829.380000 149.255000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.38 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 93.040000 829.380000 93.340000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.221 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.62 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 828.580000 37.125000 829.380000 37.425000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2047.78 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.220000 0.800000 10.520000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.273 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2048.02 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.590000 0.800000 20.890000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 379.131 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2046.66 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 201.055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1076.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.350000 0.800000 30.650000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 770.675000 368.060000 772.415000 762.840000 ;
      LAYER met4 ;
        RECT 295.355000 368.060000 297.095000 762.840000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 298.755000 371.460000 300.495000 759.440000 ;
      LAYER met4 ;
        RECT 767.275000 371.460000 769.015000 759.440000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 829.380000 820.080000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 829.380000 820.080000 ;
    LAYER met2 ;
      RECT 820.160000 819.450000 829.380000 820.080000 ;
      RECT 797.685000 819.450000 819.740000 820.080000 ;
      RECT 765.785000 819.450000 797.265000 820.080000 ;
      RECT 733.885000 819.450000 765.365000 820.080000 ;
      RECT 701.990000 819.450000 733.465000 820.080000 ;
      RECT 670.090000 819.450000 701.570000 820.080000 ;
      RECT 638.190000 819.450000 669.670000 820.080000 ;
      RECT 606.290000 819.450000 637.770000 820.080000 ;
      RECT 574.390000 819.450000 605.870000 820.080000 ;
      RECT 542.495000 819.450000 573.970000 820.080000 ;
      RECT 510.595000 819.450000 542.075000 820.080000 ;
      RECT 478.695000 819.450000 510.175000 820.080000 ;
      RECT 446.795000 819.450000 478.275000 820.080000 ;
      RECT 414.895000 819.450000 446.375000 820.080000 ;
      RECT 383.000000 819.450000 414.475000 820.080000 ;
      RECT 351.100000 819.450000 382.580000 820.080000 ;
      RECT 319.200000 819.450000 350.680000 820.080000 ;
      RECT 287.300000 819.450000 318.780000 820.080000 ;
      RECT 255.400000 819.450000 286.880000 820.080000 ;
      RECT 223.505000 819.450000 254.980000 820.080000 ;
      RECT 191.605000 819.450000 223.085000 820.080000 ;
      RECT 159.705000 819.450000 191.185000 820.080000 ;
      RECT 127.805000 819.450000 159.285000 820.080000 ;
      RECT 95.905000 819.450000 127.385000 820.080000 ;
      RECT 64.010000 819.450000 95.485000 820.080000 ;
      RECT 32.110000 819.450000 63.590000 820.080000 ;
      RECT 10.560000 819.450000 31.690000 820.080000 ;
      RECT 0.000000 819.450000 10.140000 820.080000 ;
      RECT 0.000000 10.240000 829.380000 819.450000 ;
      RECT 0.630000 9.820000 829.380000 10.240000 ;
      RECT 0.000000 0.630000 829.380000 9.820000 ;
      RECT 827.860000 0.000000 829.380000 0.630000 ;
      RECT 826.160000 0.000000 827.440000 0.630000 ;
      RECT 824.465000 0.000000 825.740000 0.630000 ;
      RECT 822.770000 0.000000 824.045000 0.630000 ;
      RECT 821.075000 0.000000 822.350000 0.630000 ;
      RECT 819.380000 0.000000 820.655000 0.630000 ;
      RECT 818.780000 0.000000 818.960000 0.630000 ;
      RECT 817.680000 0.000000 818.360000 0.630000 ;
      RECT 815.985000 0.000000 817.260000 0.630000 ;
      RECT 814.290000 0.000000 815.565000 0.630000 ;
      RECT 812.595000 0.000000 813.870000 0.630000 ;
      RECT 810.900000 0.000000 812.175000 0.630000 ;
      RECT 809.200000 0.000000 810.480000 0.630000 ;
      RECT 807.505000 0.000000 808.780000 0.630000 ;
      RECT 805.810000 0.000000 807.085000 0.630000 ;
      RECT 804.115000 0.000000 805.390000 0.630000 ;
      RECT 802.420000 0.000000 803.695000 0.630000 ;
      RECT 800.720000 0.000000 802.000000 0.630000 ;
      RECT 799.025000 0.000000 800.300000 0.630000 ;
      RECT 797.330000 0.000000 798.605000 0.630000 ;
      RECT 795.635000 0.000000 796.910000 0.630000 ;
      RECT 793.940000 0.000000 795.215000 0.630000 ;
      RECT 792.240000 0.000000 793.520000 0.630000 ;
      RECT 790.545000 0.000000 791.820000 0.630000 ;
      RECT 788.850000 0.000000 790.125000 0.630000 ;
      RECT 787.155000 0.000000 788.430000 0.630000 ;
      RECT 785.460000 0.000000 786.735000 0.630000 ;
      RECT 783.760000 0.000000 785.040000 0.630000 ;
      RECT 782.065000 0.000000 783.340000 0.630000 ;
      RECT 780.370000 0.000000 781.645000 0.630000 ;
      RECT 778.675000 0.000000 779.950000 0.630000 ;
      RECT 776.980000 0.000000 778.255000 0.630000 ;
      RECT 775.280000 0.000000 776.560000 0.630000 ;
      RECT 773.585000 0.000000 774.860000 0.630000 ;
      RECT 771.890000 0.000000 773.165000 0.630000 ;
      RECT 770.195000 0.000000 771.470000 0.630000 ;
      RECT 768.500000 0.000000 769.775000 0.630000 ;
      RECT 766.800000 0.000000 768.080000 0.630000 ;
      RECT 765.105000 0.000000 766.380000 0.630000 ;
      RECT 763.410000 0.000000 764.685000 0.630000 ;
      RECT 761.715000 0.000000 762.990000 0.630000 ;
      RECT 760.020000 0.000000 761.295000 0.630000 ;
      RECT 758.320000 0.000000 759.600000 0.630000 ;
      RECT 756.625000 0.000000 757.900000 0.630000 ;
      RECT 754.930000 0.000000 756.205000 0.630000 ;
      RECT 753.235000 0.000000 754.510000 0.630000 ;
      RECT 751.540000 0.000000 752.815000 0.630000 ;
      RECT 749.840000 0.000000 751.120000 0.630000 ;
      RECT 748.145000 0.000000 749.420000 0.630000 ;
      RECT 746.450000 0.000000 747.725000 0.630000 ;
      RECT 744.755000 0.000000 746.030000 0.630000 ;
      RECT 743.060000 0.000000 744.335000 0.630000 ;
      RECT 741.360000 0.000000 742.640000 0.630000 ;
      RECT 739.665000 0.000000 740.940000 0.630000 ;
      RECT 737.970000 0.000000 739.245000 0.630000 ;
      RECT 736.275000 0.000000 737.550000 0.630000 ;
      RECT 734.580000 0.000000 735.855000 0.630000 ;
      RECT 732.880000 0.000000 734.160000 0.630000 ;
      RECT 731.185000 0.000000 732.460000 0.630000 ;
      RECT 729.490000 0.000000 730.765000 0.630000 ;
      RECT 727.795000 0.000000 729.070000 0.630000 ;
      RECT 726.100000 0.000000 727.375000 0.630000 ;
      RECT 724.400000 0.000000 725.680000 0.630000 ;
      RECT 722.705000 0.000000 723.980000 0.630000 ;
      RECT 721.010000 0.000000 722.285000 0.630000 ;
      RECT 719.315000 0.000000 720.590000 0.630000 ;
      RECT 717.620000 0.000000 718.895000 0.630000 ;
      RECT 715.920000 0.000000 717.200000 0.630000 ;
      RECT 714.225000 0.000000 715.500000 0.630000 ;
      RECT 712.530000 0.000000 713.805000 0.630000 ;
      RECT 710.835000 0.000000 712.110000 0.630000 ;
      RECT 709.140000 0.000000 710.415000 0.630000 ;
      RECT 707.440000 0.000000 708.720000 0.630000 ;
      RECT 705.745000 0.000000 707.020000 0.630000 ;
      RECT 704.050000 0.000000 705.325000 0.630000 ;
      RECT 702.355000 0.000000 703.630000 0.630000 ;
      RECT 700.660000 0.000000 701.935000 0.630000 ;
      RECT 698.960000 0.000000 700.240000 0.630000 ;
      RECT 697.265000 0.000000 698.540000 0.630000 ;
      RECT 695.570000 0.000000 696.845000 0.630000 ;
      RECT 693.875000 0.000000 695.150000 0.630000 ;
      RECT 692.180000 0.000000 693.455000 0.630000 ;
      RECT 690.480000 0.000000 691.760000 0.630000 ;
      RECT 688.785000 0.000000 690.060000 0.630000 ;
      RECT 687.090000 0.000000 688.365000 0.630000 ;
      RECT 685.395000 0.000000 686.670000 0.630000 ;
      RECT 683.700000 0.000000 684.975000 0.630000 ;
      RECT 682.000000 0.000000 683.280000 0.630000 ;
      RECT 680.305000 0.000000 681.580000 0.630000 ;
      RECT 678.610000 0.000000 679.885000 0.630000 ;
      RECT 676.915000 0.000000 678.190000 0.630000 ;
      RECT 675.220000 0.000000 676.495000 0.630000 ;
      RECT 673.520000 0.000000 674.800000 0.630000 ;
      RECT 671.825000 0.000000 673.100000 0.630000 ;
      RECT 670.130000 0.000000 671.405000 0.630000 ;
      RECT 668.435000 0.000000 669.710000 0.630000 ;
      RECT 666.740000 0.000000 668.015000 0.630000 ;
      RECT 665.040000 0.000000 666.320000 0.630000 ;
      RECT 663.345000 0.000000 664.620000 0.630000 ;
      RECT 661.650000 0.000000 662.925000 0.630000 ;
      RECT 659.955000 0.000000 661.230000 0.630000 ;
      RECT 658.260000 0.000000 659.535000 0.630000 ;
      RECT 656.560000 0.000000 657.840000 0.630000 ;
      RECT 654.865000 0.000000 656.140000 0.630000 ;
      RECT 653.170000 0.000000 654.445000 0.630000 ;
      RECT 651.475000 0.000000 652.750000 0.630000 ;
      RECT 649.780000 0.000000 651.055000 0.630000 ;
      RECT 648.080000 0.000000 649.360000 0.630000 ;
      RECT 646.385000 0.000000 647.660000 0.630000 ;
      RECT 644.690000 0.000000 645.965000 0.630000 ;
      RECT 642.995000 0.000000 644.270000 0.630000 ;
      RECT 641.300000 0.000000 642.575000 0.630000 ;
      RECT 639.600000 0.000000 640.880000 0.630000 ;
      RECT 637.905000 0.000000 639.180000 0.630000 ;
      RECT 636.210000 0.000000 637.485000 0.630000 ;
      RECT 634.515000 0.000000 635.790000 0.630000 ;
      RECT 632.820000 0.000000 634.095000 0.630000 ;
      RECT 631.120000 0.000000 632.400000 0.630000 ;
      RECT 629.425000 0.000000 630.700000 0.630000 ;
      RECT 627.730000 0.000000 629.005000 0.630000 ;
      RECT 626.035000 0.000000 627.310000 0.630000 ;
      RECT 624.340000 0.000000 625.615000 0.630000 ;
      RECT 622.640000 0.000000 623.920000 0.630000 ;
      RECT 620.945000 0.000000 622.220000 0.630000 ;
      RECT 619.250000 0.000000 620.525000 0.630000 ;
      RECT 617.555000 0.000000 618.830000 0.630000 ;
      RECT 615.860000 0.000000 617.135000 0.630000 ;
      RECT 614.160000 0.000000 615.440000 0.630000 ;
      RECT 612.465000 0.000000 613.740000 0.630000 ;
      RECT 610.770000 0.000000 612.045000 0.630000 ;
      RECT 609.075000 0.000000 610.350000 0.630000 ;
      RECT 607.380000 0.000000 608.655000 0.630000 ;
      RECT 605.680000 0.000000 606.960000 0.630000 ;
      RECT 603.985000 0.000000 605.260000 0.630000 ;
      RECT 602.290000 0.000000 603.565000 0.630000 ;
      RECT 600.595000 0.000000 601.870000 0.630000 ;
      RECT 598.900000 0.000000 600.175000 0.630000 ;
      RECT 597.200000 0.000000 598.480000 0.630000 ;
      RECT 595.505000 0.000000 596.780000 0.630000 ;
      RECT 593.810000 0.000000 595.085000 0.630000 ;
      RECT 592.115000 0.000000 593.390000 0.630000 ;
      RECT 590.420000 0.000000 591.695000 0.630000 ;
      RECT 588.720000 0.000000 590.000000 0.630000 ;
      RECT 587.025000 0.000000 588.300000 0.630000 ;
      RECT 585.330000 0.000000 586.605000 0.630000 ;
      RECT 583.635000 0.000000 584.910000 0.630000 ;
      RECT 581.940000 0.000000 583.215000 0.630000 ;
      RECT 580.240000 0.000000 581.520000 0.630000 ;
      RECT 578.545000 0.000000 579.820000 0.630000 ;
      RECT 576.850000 0.000000 578.125000 0.630000 ;
      RECT 575.155000 0.000000 576.430000 0.630000 ;
      RECT 573.460000 0.000000 574.735000 0.630000 ;
      RECT 571.760000 0.000000 573.040000 0.630000 ;
      RECT 570.065000 0.000000 571.340000 0.630000 ;
      RECT 568.370000 0.000000 569.645000 0.630000 ;
      RECT 566.675000 0.000000 567.950000 0.630000 ;
      RECT 564.980000 0.000000 566.255000 0.630000 ;
      RECT 563.280000 0.000000 564.560000 0.630000 ;
      RECT 561.585000 0.000000 562.860000 0.630000 ;
      RECT 559.890000 0.000000 561.165000 0.630000 ;
      RECT 558.195000 0.000000 559.470000 0.630000 ;
      RECT 556.500000 0.000000 557.775000 0.630000 ;
      RECT 554.800000 0.000000 556.080000 0.630000 ;
      RECT 553.105000 0.000000 554.380000 0.630000 ;
      RECT 551.410000 0.000000 552.685000 0.630000 ;
      RECT 549.715000 0.000000 550.990000 0.630000 ;
      RECT 548.020000 0.000000 549.295000 0.630000 ;
      RECT 546.320000 0.000000 547.600000 0.630000 ;
      RECT 544.625000 0.000000 545.900000 0.630000 ;
      RECT 542.930000 0.000000 544.205000 0.630000 ;
      RECT 541.235000 0.000000 542.510000 0.630000 ;
      RECT 539.540000 0.000000 540.815000 0.630000 ;
      RECT 537.840000 0.000000 539.120000 0.630000 ;
      RECT 536.145000 0.000000 537.420000 0.630000 ;
      RECT 534.450000 0.000000 535.725000 0.630000 ;
      RECT 532.755000 0.000000 534.030000 0.630000 ;
      RECT 531.060000 0.000000 532.335000 0.630000 ;
      RECT 529.360000 0.000000 530.640000 0.630000 ;
      RECT 527.665000 0.000000 528.940000 0.630000 ;
      RECT 525.970000 0.000000 527.245000 0.630000 ;
      RECT 524.275000 0.000000 525.550000 0.630000 ;
      RECT 522.580000 0.000000 523.855000 0.630000 ;
      RECT 520.880000 0.000000 522.160000 0.630000 ;
      RECT 519.185000 0.000000 520.460000 0.630000 ;
      RECT 517.490000 0.000000 518.765000 0.630000 ;
      RECT 515.795000 0.000000 517.070000 0.630000 ;
      RECT 514.100000 0.000000 515.375000 0.630000 ;
      RECT 512.400000 0.000000 513.680000 0.630000 ;
      RECT 510.705000 0.000000 511.980000 0.630000 ;
      RECT 509.010000 0.000000 510.285000 0.630000 ;
      RECT 507.315000 0.000000 508.590000 0.630000 ;
      RECT 505.620000 0.000000 506.895000 0.630000 ;
      RECT 503.920000 0.000000 505.200000 0.630000 ;
      RECT 502.225000 0.000000 503.500000 0.630000 ;
      RECT 500.530000 0.000000 501.805000 0.630000 ;
      RECT 498.835000 0.000000 500.110000 0.630000 ;
      RECT 497.140000 0.000000 498.415000 0.630000 ;
      RECT 495.440000 0.000000 496.720000 0.630000 ;
      RECT 493.745000 0.000000 495.020000 0.630000 ;
      RECT 492.050000 0.000000 493.325000 0.630000 ;
      RECT 490.355000 0.000000 491.630000 0.630000 ;
      RECT 488.660000 0.000000 489.935000 0.630000 ;
      RECT 486.960000 0.000000 488.240000 0.630000 ;
      RECT 485.265000 0.000000 486.540000 0.630000 ;
      RECT 483.570000 0.000000 484.845000 0.630000 ;
      RECT 481.875000 0.000000 483.150000 0.630000 ;
      RECT 480.180000 0.000000 481.455000 0.630000 ;
      RECT 478.480000 0.000000 479.760000 0.630000 ;
      RECT 476.785000 0.000000 478.060000 0.630000 ;
      RECT 475.090000 0.000000 476.365000 0.630000 ;
      RECT 473.395000 0.000000 474.670000 0.630000 ;
      RECT 471.700000 0.000000 472.975000 0.630000 ;
      RECT 470.000000 0.000000 471.280000 0.630000 ;
      RECT 468.305000 0.000000 469.580000 0.630000 ;
      RECT 466.610000 0.000000 467.885000 0.630000 ;
      RECT 464.915000 0.000000 466.190000 0.630000 ;
      RECT 463.220000 0.000000 464.495000 0.630000 ;
      RECT 461.520000 0.000000 462.800000 0.630000 ;
      RECT 459.825000 0.000000 461.100000 0.630000 ;
      RECT 458.130000 0.000000 459.405000 0.630000 ;
      RECT 456.435000 0.000000 457.710000 0.630000 ;
      RECT 454.740000 0.000000 456.015000 0.630000 ;
      RECT 453.040000 0.000000 454.320000 0.630000 ;
      RECT 451.345000 0.000000 452.620000 0.630000 ;
      RECT 449.650000 0.000000 450.925000 0.630000 ;
      RECT 447.955000 0.000000 449.230000 0.630000 ;
      RECT 446.260000 0.000000 447.535000 0.630000 ;
      RECT 444.560000 0.000000 445.840000 0.630000 ;
      RECT 442.865000 0.000000 444.140000 0.630000 ;
      RECT 441.170000 0.000000 442.445000 0.630000 ;
      RECT 439.475000 0.000000 440.750000 0.630000 ;
      RECT 437.780000 0.000000 439.055000 0.630000 ;
      RECT 436.080000 0.000000 437.360000 0.630000 ;
      RECT 434.385000 0.000000 435.660000 0.630000 ;
      RECT 432.690000 0.000000 433.965000 0.630000 ;
      RECT 430.995000 0.000000 432.270000 0.630000 ;
      RECT 429.300000 0.000000 430.575000 0.630000 ;
      RECT 427.600000 0.000000 428.880000 0.630000 ;
      RECT 425.905000 0.000000 427.180000 0.630000 ;
      RECT 424.210000 0.000000 425.485000 0.630000 ;
      RECT 422.515000 0.000000 423.790000 0.630000 ;
      RECT 420.820000 0.000000 422.095000 0.630000 ;
      RECT 419.120000 0.000000 420.400000 0.630000 ;
      RECT 417.425000 0.000000 418.700000 0.630000 ;
      RECT 415.730000 0.000000 417.005000 0.630000 ;
      RECT 414.035000 0.000000 415.310000 0.630000 ;
      RECT 412.340000 0.000000 413.615000 0.630000 ;
      RECT 410.640000 0.000000 411.920000 0.630000 ;
      RECT 408.945000 0.000000 410.220000 0.630000 ;
      RECT 407.250000 0.000000 408.525000 0.630000 ;
      RECT 405.555000 0.000000 406.830000 0.630000 ;
      RECT 403.860000 0.000000 405.135000 0.630000 ;
      RECT 402.160000 0.000000 403.440000 0.630000 ;
      RECT 400.465000 0.000000 401.740000 0.630000 ;
      RECT 398.770000 0.000000 400.045000 0.630000 ;
      RECT 397.075000 0.000000 398.350000 0.630000 ;
      RECT 395.380000 0.000000 396.655000 0.630000 ;
      RECT 393.680000 0.000000 394.960000 0.630000 ;
      RECT 391.985000 0.000000 393.260000 0.630000 ;
      RECT 390.290000 0.000000 391.565000 0.630000 ;
      RECT 388.595000 0.000000 389.870000 0.630000 ;
      RECT 386.900000 0.000000 388.175000 0.630000 ;
      RECT 385.200000 0.000000 386.480000 0.630000 ;
      RECT 383.505000 0.000000 384.780000 0.630000 ;
      RECT 381.810000 0.000000 383.085000 0.630000 ;
      RECT 380.115000 0.000000 381.390000 0.630000 ;
      RECT 378.420000 0.000000 379.695000 0.630000 ;
      RECT 376.720000 0.000000 378.000000 0.630000 ;
      RECT 375.025000 0.000000 376.300000 0.630000 ;
      RECT 373.330000 0.000000 374.605000 0.630000 ;
      RECT 371.635000 0.000000 372.910000 0.630000 ;
      RECT 369.940000 0.000000 371.215000 0.630000 ;
      RECT 368.240000 0.000000 369.520000 0.630000 ;
      RECT 366.545000 0.000000 367.820000 0.630000 ;
      RECT 364.850000 0.000000 366.125000 0.630000 ;
      RECT 363.155000 0.000000 364.430000 0.630000 ;
      RECT 361.460000 0.000000 362.735000 0.630000 ;
      RECT 359.760000 0.000000 361.040000 0.630000 ;
      RECT 358.065000 0.000000 359.340000 0.630000 ;
      RECT 356.370000 0.000000 357.645000 0.630000 ;
      RECT 354.675000 0.000000 355.950000 0.630000 ;
      RECT 352.980000 0.000000 354.255000 0.630000 ;
      RECT 351.280000 0.000000 352.560000 0.630000 ;
      RECT 349.585000 0.000000 350.860000 0.630000 ;
      RECT 347.890000 0.000000 349.165000 0.630000 ;
      RECT 346.195000 0.000000 347.470000 0.630000 ;
      RECT 344.500000 0.000000 345.775000 0.630000 ;
      RECT 342.800000 0.000000 344.080000 0.630000 ;
      RECT 341.105000 0.000000 342.380000 0.630000 ;
      RECT 339.410000 0.000000 340.685000 0.630000 ;
      RECT 337.715000 0.000000 338.990000 0.630000 ;
      RECT 336.020000 0.000000 337.295000 0.630000 ;
      RECT 334.320000 0.000000 335.600000 0.630000 ;
      RECT 332.625000 0.000000 333.900000 0.630000 ;
      RECT 330.930000 0.000000 332.205000 0.630000 ;
      RECT 329.235000 0.000000 330.510000 0.630000 ;
      RECT 327.540000 0.000000 328.815000 0.630000 ;
      RECT 325.840000 0.000000 327.120000 0.630000 ;
      RECT 324.145000 0.000000 325.420000 0.630000 ;
      RECT 322.450000 0.000000 323.725000 0.630000 ;
      RECT 320.755000 0.000000 322.030000 0.630000 ;
      RECT 319.060000 0.000000 320.335000 0.630000 ;
      RECT 317.360000 0.000000 318.640000 0.630000 ;
      RECT 315.665000 0.000000 316.940000 0.630000 ;
      RECT 313.970000 0.000000 315.245000 0.630000 ;
      RECT 312.275000 0.000000 313.550000 0.630000 ;
      RECT 310.580000 0.000000 311.855000 0.630000 ;
      RECT 308.880000 0.000000 310.160000 0.630000 ;
      RECT 307.185000 0.000000 308.460000 0.630000 ;
      RECT 305.490000 0.000000 306.765000 0.630000 ;
      RECT 303.795000 0.000000 305.070000 0.630000 ;
      RECT 302.100000 0.000000 303.375000 0.630000 ;
      RECT 300.400000 0.000000 301.680000 0.630000 ;
      RECT 298.705000 0.000000 299.980000 0.630000 ;
      RECT 297.010000 0.000000 298.285000 0.630000 ;
      RECT 295.315000 0.000000 296.590000 0.630000 ;
      RECT 293.620000 0.000000 294.895000 0.630000 ;
      RECT 291.920000 0.000000 293.200000 0.630000 ;
      RECT 290.225000 0.000000 291.500000 0.630000 ;
      RECT 288.530000 0.000000 289.805000 0.630000 ;
      RECT 286.835000 0.000000 288.110000 0.630000 ;
      RECT 285.140000 0.000000 286.415000 0.630000 ;
      RECT 283.440000 0.000000 284.720000 0.630000 ;
      RECT 281.745000 0.000000 283.020000 0.630000 ;
      RECT 280.050000 0.000000 281.325000 0.630000 ;
      RECT 278.355000 0.000000 279.630000 0.630000 ;
      RECT 276.660000 0.000000 277.935000 0.630000 ;
      RECT 274.960000 0.000000 276.240000 0.630000 ;
      RECT 273.265000 0.000000 274.540000 0.630000 ;
      RECT 271.570000 0.000000 272.845000 0.630000 ;
      RECT 269.875000 0.000000 271.150000 0.630000 ;
      RECT 268.180000 0.000000 269.455000 0.630000 ;
      RECT 266.480000 0.000000 267.760000 0.630000 ;
      RECT 264.785000 0.000000 266.060000 0.630000 ;
      RECT 263.090000 0.000000 264.365000 0.630000 ;
      RECT 261.395000 0.000000 262.670000 0.630000 ;
      RECT 259.700000 0.000000 260.975000 0.630000 ;
      RECT 258.000000 0.000000 259.280000 0.630000 ;
      RECT 256.305000 0.000000 257.580000 0.630000 ;
      RECT 254.610000 0.000000 255.885000 0.630000 ;
      RECT 252.915000 0.000000 254.190000 0.630000 ;
      RECT 251.220000 0.000000 252.495000 0.630000 ;
      RECT 249.520000 0.000000 250.800000 0.630000 ;
      RECT 247.825000 0.000000 249.100000 0.630000 ;
      RECT 246.130000 0.000000 247.405000 0.630000 ;
      RECT 244.435000 0.000000 245.710000 0.630000 ;
      RECT 242.740000 0.000000 244.015000 0.630000 ;
      RECT 241.040000 0.000000 242.320000 0.630000 ;
      RECT 239.345000 0.000000 240.620000 0.630000 ;
      RECT 237.650000 0.000000 238.925000 0.630000 ;
      RECT 235.955000 0.000000 237.230000 0.630000 ;
      RECT 234.260000 0.000000 235.535000 0.630000 ;
      RECT 232.560000 0.000000 233.840000 0.630000 ;
      RECT 230.865000 0.000000 232.140000 0.630000 ;
      RECT 229.170000 0.000000 230.445000 0.630000 ;
      RECT 227.475000 0.000000 228.750000 0.630000 ;
      RECT 225.780000 0.000000 227.055000 0.630000 ;
      RECT 224.080000 0.000000 225.360000 0.630000 ;
      RECT 222.385000 0.000000 223.660000 0.630000 ;
      RECT 220.690000 0.000000 221.965000 0.630000 ;
      RECT 218.995000 0.000000 220.270000 0.630000 ;
      RECT 217.300000 0.000000 218.575000 0.630000 ;
      RECT 215.600000 0.000000 216.880000 0.630000 ;
      RECT 213.905000 0.000000 215.180000 0.630000 ;
      RECT 212.210000 0.000000 213.485000 0.630000 ;
      RECT 210.515000 0.000000 211.790000 0.630000 ;
      RECT 208.820000 0.000000 210.095000 0.630000 ;
      RECT 207.120000 0.000000 208.400000 0.630000 ;
      RECT 205.425000 0.000000 206.700000 0.630000 ;
      RECT 203.730000 0.000000 205.005000 0.630000 ;
      RECT 202.035000 0.000000 203.310000 0.630000 ;
      RECT 200.340000 0.000000 201.615000 0.630000 ;
      RECT 198.640000 0.000000 199.920000 0.630000 ;
      RECT 196.945000 0.000000 198.220000 0.630000 ;
      RECT 195.250000 0.000000 196.525000 0.630000 ;
      RECT 193.555000 0.000000 194.830000 0.630000 ;
      RECT 191.860000 0.000000 193.135000 0.630000 ;
      RECT 190.160000 0.000000 191.440000 0.630000 ;
      RECT 188.465000 0.000000 189.740000 0.630000 ;
      RECT 186.770000 0.000000 188.045000 0.630000 ;
      RECT 185.075000 0.000000 186.350000 0.630000 ;
      RECT 183.380000 0.000000 184.655000 0.630000 ;
      RECT 181.680000 0.000000 182.960000 0.630000 ;
      RECT 179.985000 0.000000 181.260000 0.630000 ;
      RECT 178.290000 0.000000 179.565000 0.630000 ;
      RECT 176.595000 0.000000 177.870000 0.630000 ;
      RECT 174.900000 0.000000 176.175000 0.630000 ;
      RECT 173.200000 0.000000 174.480000 0.630000 ;
      RECT 171.505000 0.000000 172.780000 0.630000 ;
      RECT 169.810000 0.000000 171.085000 0.630000 ;
      RECT 168.115000 0.000000 169.390000 0.630000 ;
      RECT 166.420000 0.000000 167.695000 0.630000 ;
      RECT 164.720000 0.000000 166.000000 0.630000 ;
      RECT 163.025000 0.000000 164.300000 0.630000 ;
      RECT 161.330000 0.000000 162.605000 0.630000 ;
      RECT 159.635000 0.000000 160.910000 0.630000 ;
      RECT 157.940000 0.000000 159.215000 0.630000 ;
      RECT 156.240000 0.000000 157.520000 0.630000 ;
      RECT 154.545000 0.000000 155.820000 0.630000 ;
      RECT 152.850000 0.000000 154.125000 0.630000 ;
      RECT 151.155000 0.000000 152.430000 0.630000 ;
      RECT 149.460000 0.000000 150.735000 0.630000 ;
      RECT 147.760000 0.000000 149.040000 0.630000 ;
      RECT 146.065000 0.000000 147.340000 0.630000 ;
      RECT 144.370000 0.000000 145.645000 0.630000 ;
      RECT 142.675000 0.000000 143.950000 0.630000 ;
      RECT 140.980000 0.000000 142.255000 0.630000 ;
      RECT 139.280000 0.000000 140.560000 0.630000 ;
      RECT 137.585000 0.000000 138.860000 0.630000 ;
      RECT 135.890000 0.000000 137.165000 0.630000 ;
      RECT 134.195000 0.000000 135.470000 0.630000 ;
      RECT 132.500000 0.000000 133.775000 0.630000 ;
      RECT 130.800000 0.000000 132.080000 0.630000 ;
      RECT 129.105000 0.000000 130.380000 0.630000 ;
      RECT 127.410000 0.000000 128.685000 0.630000 ;
      RECT 125.715000 0.000000 126.990000 0.630000 ;
      RECT 124.020000 0.000000 125.295000 0.630000 ;
      RECT 122.320000 0.000000 123.600000 0.630000 ;
      RECT 120.625000 0.000000 121.900000 0.630000 ;
      RECT 118.930000 0.000000 120.205000 0.630000 ;
      RECT 117.235000 0.000000 118.510000 0.630000 ;
      RECT 115.540000 0.000000 116.815000 0.630000 ;
      RECT 113.840000 0.000000 115.120000 0.630000 ;
      RECT 112.145000 0.000000 113.420000 0.630000 ;
      RECT 110.450000 0.000000 111.725000 0.630000 ;
      RECT 108.755000 0.000000 110.030000 0.630000 ;
      RECT 107.060000 0.000000 108.335000 0.630000 ;
      RECT 105.360000 0.000000 106.640000 0.630000 ;
      RECT 103.665000 0.000000 104.940000 0.630000 ;
      RECT 101.970000 0.000000 103.245000 0.630000 ;
      RECT 100.275000 0.000000 101.550000 0.630000 ;
      RECT 98.580000 0.000000 99.855000 0.630000 ;
      RECT 96.880000 0.000000 98.160000 0.630000 ;
      RECT 95.185000 0.000000 96.460000 0.630000 ;
      RECT 93.490000 0.000000 94.765000 0.630000 ;
      RECT 91.795000 0.000000 93.070000 0.630000 ;
      RECT 90.100000 0.000000 91.375000 0.630000 ;
      RECT 88.400000 0.000000 89.680000 0.630000 ;
      RECT 86.705000 0.000000 87.980000 0.630000 ;
      RECT 85.010000 0.000000 86.285000 0.630000 ;
      RECT 83.315000 0.000000 84.590000 0.630000 ;
      RECT 81.620000 0.000000 82.895000 0.630000 ;
      RECT 79.920000 0.000000 81.200000 0.630000 ;
      RECT 78.225000 0.000000 79.500000 0.630000 ;
      RECT 76.530000 0.000000 77.805000 0.630000 ;
      RECT 74.835000 0.000000 76.110000 0.630000 ;
      RECT 73.140000 0.000000 74.415000 0.630000 ;
      RECT 71.440000 0.000000 72.720000 0.630000 ;
      RECT 69.745000 0.000000 71.020000 0.630000 ;
      RECT 68.050000 0.000000 69.325000 0.630000 ;
      RECT 66.355000 0.000000 67.630000 0.630000 ;
      RECT 64.660000 0.000000 65.935000 0.630000 ;
      RECT 62.960000 0.000000 64.240000 0.630000 ;
      RECT 61.265000 0.000000 62.540000 0.630000 ;
      RECT 59.570000 0.000000 60.845000 0.630000 ;
      RECT 57.875000 0.000000 59.150000 0.630000 ;
      RECT 56.180000 0.000000 57.455000 0.630000 ;
      RECT 54.480000 0.000000 55.760000 0.630000 ;
      RECT 52.785000 0.000000 54.060000 0.630000 ;
      RECT 51.090000 0.000000 52.365000 0.630000 ;
      RECT 49.395000 0.000000 50.670000 0.630000 ;
      RECT 47.700000 0.000000 48.975000 0.630000 ;
      RECT 46.000000 0.000000 47.280000 0.630000 ;
      RECT 44.305000 0.000000 45.580000 0.630000 ;
      RECT 42.610000 0.000000 43.885000 0.630000 ;
      RECT 40.915000 0.000000 42.190000 0.630000 ;
      RECT 39.220000 0.000000 40.495000 0.630000 ;
      RECT 37.520000 0.000000 38.800000 0.630000 ;
      RECT 35.825000 0.000000 37.100000 0.630000 ;
      RECT 34.130000 0.000000 35.405000 0.630000 ;
      RECT 32.435000 0.000000 33.710000 0.630000 ;
      RECT 30.740000 0.000000 32.015000 0.630000 ;
      RECT 29.040000 0.000000 30.320000 0.630000 ;
      RECT 27.345000 0.000000 28.620000 0.630000 ;
      RECT 25.650000 0.000000 26.925000 0.630000 ;
      RECT 23.955000 0.000000 25.230000 0.630000 ;
      RECT 22.260000 0.000000 23.535000 0.630000 ;
      RECT 20.560000 0.000000 21.840000 0.630000 ;
      RECT 18.865000 0.000000 20.140000 0.630000 ;
      RECT 17.170000 0.000000 18.445000 0.630000 ;
      RECT 15.475000 0.000000 16.750000 0.630000 ;
      RECT 13.780000 0.000000 15.055000 0.630000 ;
      RECT 12.080000 0.000000 13.360000 0.630000 ;
      RECT 10.385000 0.000000 11.660000 0.630000 ;
      RECT 8.690000 0.000000 9.965000 0.630000 ;
      RECT 6.995000 0.000000 8.270000 0.630000 ;
      RECT 5.300000 0.000000 6.575000 0.630000 ;
      RECT 3.600000 0.000000 4.880000 0.630000 ;
      RECT 1.905000 0.000000 3.180000 0.630000 ;
      RECT 0.000000 0.000000 1.485000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 819.390000 828.280000 820.080000 ;
      RECT 0.000000 801.885000 829.380000 819.390000 ;
      RECT 0.000000 800.985000 828.280000 801.885000 ;
      RECT 0.000000 800.490000 829.380000 800.985000 ;
      RECT 1.100000 799.590000 829.380000 800.490000 ;
      RECT 0.000000 783.245000 829.380000 799.590000 ;
      RECT 0.000000 782.345000 828.280000 783.245000 ;
      RECT 0.000000 780.490000 829.380000 782.345000 ;
      RECT 1.100000 779.590000 829.380000 780.490000 ;
      RECT 0.000000 764.610000 829.380000 779.590000 ;
      RECT 0.000000 763.710000 828.280000 764.610000 ;
      RECT 0.000000 760.490000 829.380000 763.710000 ;
      RECT 1.100000 759.590000 829.380000 760.490000 ;
      RECT 0.000000 745.970000 829.380000 759.590000 ;
      RECT 0.000000 745.070000 828.280000 745.970000 ;
      RECT 0.000000 740.485000 829.380000 745.070000 ;
      RECT 1.100000 739.585000 829.380000 740.485000 ;
      RECT 0.000000 727.330000 829.380000 739.585000 ;
      RECT 0.000000 726.430000 828.280000 727.330000 ;
      RECT 0.000000 720.485000 829.380000 726.430000 ;
      RECT 1.100000 719.585000 829.380000 720.485000 ;
      RECT 0.000000 708.695000 829.380000 719.585000 ;
      RECT 0.000000 707.795000 828.280000 708.695000 ;
      RECT 0.000000 700.485000 829.380000 707.795000 ;
      RECT 1.100000 699.585000 829.380000 700.485000 ;
      RECT 0.000000 690.055000 829.380000 699.585000 ;
      RECT 0.000000 689.155000 828.280000 690.055000 ;
      RECT 0.000000 680.485000 829.380000 689.155000 ;
      RECT 1.100000 679.585000 829.380000 680.485000 ;
      RECT 0.000000 671.420000 829.380000 679.585000 ;
      RECT 0.000000 670.520000 828.280000 671.420000 ;
      RECT 0.000000 660.485000 829.380000 670.520000 ;
      RECT 1.100000 659.585000 829.380000 660.485000 ;
      RECT 0.000000 652.780000 829.380000 659.585000 ;
      RECT 0.000000 651.880000 828.280000 652.780000 ;
      RECT 0.000000 640.480000 829.380000 651.880000 ;
      RECT 1.100000 639.580000 829.380000 640.480000 ;
      RECT 0.000000 634.140000 829.380000 639.580000 ;
      RECT 0.000000 633.240000 828.280000 634.140000 ;
      RECT 0.000000 620.480000 829.380000 633.240000 ;
      RECT 1.100000 619.580000 829.380000 620.480000 ;
      RECT 0.000000 615.505000 829.380000 619.580000 ;
      RECT 0.000000 614.605000 828.280000 615.505000 ;
      RECT 0.000000 600.480000 829.380000 614.605000 ;
      RECT 1.100000 599.580000 829.380000 600.480000 ;
      RECT 0.000000 596.865000 829.380000 599.580000 ;
      RECT 0.000000 595.965000 828.280000 596.865000 ;
      RECT 0.000000 580.480000 829.380000 595.965000 ;
      RECT 1.100000 579.580000 829.380000 580.480000 ;
      RECT 0.000000 578.230000 829.380000 579.580000 ;
      RECT 0.000000 577.330000 828.280000 578.230000 ;
      RECT 0.000000 560.480000 829.380000 577.330000 ;
      RECT 1.100000 559.590000 829.380000 560.480000 ;
      RECT 1.100000 559.580000 828.280000 559.590000 ;
      RECT 0.000000 558.690000 828.280000 559.580000 ;
      RECT 0.000000 540.950000 829.380000 558.690000 ;
      RECT 0.000000 540.475000 828.280000 540.950000 ;
      RECT 1.100000 540.050000 828.280000 540.475000 ;
      RECT 1.100000 539.575000 829.380000 540.050000 ;
      RECT 0.000000 522.315000 829.380000 539.575000 ;
      RECT 0.000000 521.415000 828.280000 522.315000 ;
      RECT 0.000000 520.475000 829.380000 521.415000 ;
      RECT 1.100000 519.575000 829.380000 520.475000 ;
      RECT 0.000000 503.675000 829.380000 519.575000 ;
      RECT 0.000000 502.775000 828.280000 503.675000 ;
      RECT 0.000000 500.475000 829.380000 502.775000 ;
      RECT 1.100000 499.575000 829.380000 500.475000 ;
      RECT 0.000000 485.040000 829.380000 499.575000 ;
      RECT 0.000000 484.140000 828.280000 485.040000 ;
      RECT 0.000000 480.475000 829.380000 484.140000 ;
      RECT 1.100000 479.575000 829.380000 480.475000 ;
      RECT 0.000000 466.400000 829.380000 479.575000 ;
      RECT 0.000000 465.500000 828.280000 466.400000 ;
      RECT 0.000000 460.475000 829.380000 465.500000 ;
      RECT 1.100000 459.575000 829.380000 460.475000 ;
      RECT 0.000000 447.760000 829.380000 459.575000 ;
      RECT 0.000000 446.860000 828.280000 447.760000 ;
      RECT 0.000000 440.470000 829.380000 446.860000 ;
      RECT 1.100000 439.570000 829.380000 440.470000 ;
      RECT 0.000000 429.125000 829.380000 439.570000 ;
      RECT 0.000000 428.225000 828.280000 429.125000 ;
      RECT 0.000000 420.470000 829.380000 428.225000 ;
      RECT 1.100000 419.570000 829.380000 420.470000 ;
      RECT 0.000000 410.485000 829.380000 419.570000 ;
      RECT 0.000000 409.585000 828.280000 410.485000 ;
      RECT 0.000000 400.470000 829.380000 409.585000 ;
      RECT 1.100000 399.570000 829.380000 400.470000 ;
      RECT 0.000000 391.850000 829.380000 399.570000 ;
      RECT 0.000000 390.950000 828.280000 391.850000 ;
      RECT 0.000000 380.470000 829.380000 390.950000 ;
      RECT 1.100000 379.570000 829.380000 380.470000 ;
      RECT 0.000000 373.210000 829.380000 379.570000 ;
      RECT 0.000000 372.310000 828.280000 373.210000 ;
      RECT 0.000000 360.470000 829.380000 372.310000 ;
      RECT 1.100000 359.570000 829.380000 360.470000 ;
      RECT 0.000000 354.570000 829.380000 359.570000 ;
      RECT 0.000000 353.670000 828.280000 354.570000 ;
      RECT 0.000000 340.465000 829.380000 353.670000 ;
      RECT 1.100000 339.565000 829.380000 340.465000 ;
      RECT 0.000000 335.935000 829.380000 339.565000 ;
      RECT 0.000000 335.035000 828.280000 335.935000 ;
      RECT 0.000000 320.465000 829.380000 335.035000 ;
      RECT 1.100000 319.565000 829.380000 320.465000 ;
      RECT 0.000000 317.295000 829.380000 319.565000 ;
      RECT 0.000000 316.395000 828.280000 317.295000 ;
      RECT 0.000000 300.465000 829.380000 316.395000 ;
      RECT 1.100000 299.565000 829.380000 300.465000 ;
      RECT 0.000000 298.660000 829.380000 299.565000 ;
      RECT 0.000000 297.760000 828.280000 298.660000 ;
      RECT 0.000000 280.465000 829.380000 297.760000 ;
      RECT 1.100000 280.020000 829.380000 280.465000 ;
      RECT 1.100000 279.565000 828.280000 280.020000 ;
      RECT 0.000000 279.120000 828.280000 279.565000 ;
      RECT 0.000000 261.380000 829.380000 279.120000 ;
      RECT 0.000000 260.480000 828.280000 261.380000 ;
      RECT 0.000000 260.465000 829.380000 260.480000 ;
      RECT 1.100000 259.565000 829.380000 260.465000 ;
      RECT 0.000000 242.745000 829.380000 259.565000 ;
      RECT 0.000000 241.845000 828.280000 242.745000 ;
      RECT 0.000000 240.460000 829.380000 241.845000 ;
      RECT 1.100000 239.560000 829.380000 240.460000 ;
      RECT 0.000000 224.105000 829.380000 239.560000 ;
      RECT 0.000000 223.205000 828.280000 224.105000 ;
      RECT 0.000000 220.460000 829.380000 223.205000 ;
      RECT 1.100000 219.560000 829.380000 220.460000 ;
      RECT 0.000000 205.470000 829.380000 219.560000 ;
      RECT 0.000000 204.570000 828.280000 205.470000 ;
      RECT 0.000000 200.460000 829.380000 204.570000 ;
      RECT 1.100000 199.560000 829.380000 200.460000 ;
      RECT 0.000000 186.830000 829.380000 199.560000 ;
      RECT 0.000000 185.930000 828.280000 186.830000 ;
      RECT 0.000000 180.460000 829.380000 185.930000 ;
      RECT 1.100000 179.560000 829.380000 180.460000 ;
      RECT 0.000000 168.190000 829.380000 179.560000 ;
      RECT 0.000000 167.290000 828.280000 168.190000 ;
      RECT 0.000000 160.460000 829.380000 167.290000 ;
      RECT 1.100000 159.560000 829.380000 160.460000 ;
      RECT 0.000000 149.555000 829.380000 159.560000 ;
      RECT 0.000000 148.655000 828.280000 149.555000 ;
      RECT 0.000000 140.455000 829.380000 148.655000 ;
      RECT 1.100000 139.555000 829.380000 140.455000 ;
      RECT 0.000000 130.915000 829.380000 139.555000 ;
      RECT 0.000000 130.015000 828.280000 130.915000 ;
      RECT 0.000000 120.455000 829.380000 130.015000 ;
      RECT 1.100000 119.555000 829.380000 120.455000 ;
      RECT 0.000000 112.280000 829.380000 119.555000 ;
      RECT 0.000000 111.380000 828.280000 112.280000 ;
      RECT 0.000000 100.455000 829.380000 111.380000 ;
      RECT 1.100000 99.555000 829.380000 100.455000 ;
      RECT 0.000000 93.640000 829.380000 99.555000 ;
      RECT 0.000000 92.740000 828.280000 93.640000 ;
      RECT 0.000000 80.455000 829.380000 92.740000 ;
      RECT 1.100000 79.555000 829.380000 80.455000 ;
      RECT 0.000000 75.000000 829.380000 79.555000 ;
      RECT 0.000000 74.100000 828.280000 75.000000 ;
      RECT 0.000000 60.455000 829.380000 74.100000 ;
      RECT 1.100000 59.555000 829.380000 60.455000 ;
      RECT 0.000000 56.365000 829.380000 59.555000 ;
      RECT 0.000000 55.465000 828.280000 56.365000 ;
      RECT 0.000000 40.450000 829.380000 55.465000 ;
      RECT 1.100000 39.550000 829.380000 40.450000 ;
      RECT 0.000000 37.725000 829.380000 39.550000 ;
      RECT 0.000000 36.825000 828.280000 37.725000 ;
      RECT 0.000000 30.950000 829.380000 36.825000 ;
      RECT 1.100000 30.050000 829.380000 30.950000 ;
      RECT 0.000000 21.190000 829.380000 30.050000 ;
      RECT 1.100000 19.550000 829.380000 21.190000 ;
      RECT 0.000000 19.090000 829.380000 19.550000 ;
      RECT 0.000000 18.190000 828.280000 19.090000 ;
      RECT 0.000000 11.430000 829.380000 18.190000 ;
      RECT 1.100000 10.210000 829.380000 11.430000 ;
      RECT 1.100000 9.920000 828.280000 10.210000 ;
      RECT 0.000000 9.310000 828.280000 9.920000 ;
      RECT 0.000000 1.100000 829.380000 9.310000 ;
      RECT 10.800000 0.000000 829.380000 1.100000 ;
      RECT 0.000000 0.000000 9.900000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 0.000000 829.380000 820.080000 ;
  END
END user_proj_example

END LIBRARY
